.include ./data/sky130.sp
*For NOR2x2 --> 2 inputs, size 2 // size of each pmos cell will be 4kp, while size of nmos cell will be 2
*Instance of the cmos/pmos (source gate drain source sky130_fd_pr__esd_nfet_01v8__tt W=// L=//  )
* d g s b
*b pmos vdd
*b nmos gnd
X1 n1 a vdd vdd sky130_fd_pr__pfet_01v8 W=4000000u L=150000u
X2 c b n1 n1 sky130_fd_pr__pfet_01v8 W=4000000u L=150000u

X3 c a gnd gnd sky130_fd_pr__nfet_01v8 W=840000u L=150000u
X4 c b gnd gnd sky130_fd_pr__nfet_01v8 W=840000u L=150000u

*v(a)=0, v(b)=0, v(c)=1 correct
*v(a)=0, v(b)=1, v(c)=0 correct
*v(a)=1, v(b)=0, v(c)=0 correct
*v(a)=1, v(b)=1, v(c)=0 correct

vdd vdd gnd 1.8v
vina a gnd PULSE 1.8 0 0ps 0ps 0ps 20ns 100ns 
vinb b gnd PULSE 1.8 0 0ps 0ps 0ps 20ns 100ns

CL1 c gnd 15ff

.tran 10ps 100ns
.control
 run
 set color0=white
 set color1=black
 set xbrushwidth=2
 plot v(a), v(b), v(c)
 meas tran tpdr 
    + TRIG v(a) VAL=0.9 FALL=1
    + TARG v(c) VAL=0.9 RISE=1
 meas tran tpdf 
    + TRIG v(a) VAL=0.9 RISE=1
    + TARG v(c) VAL=0.9 FALL=1
.endc